/*******************************************************
 * Copyright (C) 2022 National Research University of Electronic Technology (MIET),
 * Institute of Microdevices and Control Systems.
 * All Rights Reserved.
 *
 * This file is part of  miriscv core.
 *
 *
 *******************************************************/

package  miriscv_cu_pkg;

  parameter NO_BYPASS = 2'd0;
  parameter BYPASS_E  = 2'd1;
  parameter BYPASS_M  = 2'd2;
  parameter BYPASS_W  = 2'd3;


endpackage :  miriscv_cu_pkg